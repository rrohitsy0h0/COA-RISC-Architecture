module Arithmetic (
    input [31:0] x,
    input [31:0] y,
    output [31:0] A_out
);
    
    f

endmodule